`define PORT_NUB_TOTAL 4
`define DATA_WIDTH 32
`define PRI_NUM_TOTAL 8
`define CRC32_LENGTH 16
`define DATABUF_HIGH_NUM 9
