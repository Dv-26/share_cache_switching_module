//端口数量
`define PORT_NUB_TOTAL 4
//数据位宽
`define DATA_WIDTH 32
//SRAM深度
`define DEPTH   1024
//数据包最大长度
`define DATA_LENGTH_MAX   256
//优先级数量
`define PRIORITY    8
`define PRI_NUM_TOTAL 8
//组合逻辑流水线优化
`define PIPELINE   1
//crc校验宽度
`define CRC32_LENGTH 16
