`define PORT_NUB_TOTAL 8
`define DATA_WIDTH 1