//端口数
`define PORT_NUB_TOTAL 4
//数据位宽
`define DATA_WIDTH 32
//SRAM深度
`define DEPTH   256
//最大包长
`define DATA_LENGTH_MAX   256
//优先级数量
`define PRIORITY    8
//是否开启流水线
`define PIPELINE   1
