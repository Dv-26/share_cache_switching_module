//端口数
`define PORT_NUB_TOTAL 4
//数据位宽
`define DATA_WIDTH 32
//SRAM深度
`define DEPTH   256
//最大包长
`define DATA_LENGTH_MAX   256
//优先级数量
`define PRIORITY    8
`define PRI_NUM_TOTAL 8
//是否开启流水线
`define PIPELINE   1
//校验码长度
`define CRC32_LENGTH 16
//包长所占位宽
`define DATABUF_HIGH_NUM 9
