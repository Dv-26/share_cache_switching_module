`ifndef SIM
    `define PORT_NUB_TOTAL 4
    `define DATA_WIDTH 6
`else
    `define PORT_NUB_TOTAL 4
    `define DATA_WIDTH 6
`endif
