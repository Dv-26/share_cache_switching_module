`define PORT_NUB_TOTAL 16
`define INPUT_DATA_WIDTH 64
`define OUTPUT_DATA_WIDTH 73
`define PRI_NUM 8
`define DATABUF_HIGH_LIMIT_NUM 256
`define CRC32_LENGTH_WIDTH 32
`define INPUT_HIGH_LIMIT_NUM 128
`define INPUT_LOW_LIMIT_NUM 8