`define PORT_NUB_TOTAL 16
`define DATA_WIDTH 1
