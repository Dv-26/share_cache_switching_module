`define PORT_NUB_TOTAL 4
`define DATA_WIDTH 1
