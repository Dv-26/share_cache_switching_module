//端口�?
`define PORT_NUB_TOTAL 8
//数据位宽
`define DATA_WIDTH 32
//SRAM深度
`define DEPTH   256
//�?大包�?
`define DATA_LENGTH_MAX   256
//优先级数�?
`define PRIORITY    8
`define PRI_NUM_TOTAL 8
//是否�?启流水线
`define PIPELINE   1
//校验码长�?
`define CRC32_LENGTH 16
//包长�?占位�?
`define DATABUF_HIGH_NUM 9
